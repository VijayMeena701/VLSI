`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:43:43 11/15/2020 
// Design Name: 
// Module Name:    array_mult 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module array_mult(
    input [15:0]c,
    input [15:0]d,
    input cin,
    output [15:0]s,
    output cout
    );


endmodule
